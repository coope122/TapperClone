module Tapper() begin
	